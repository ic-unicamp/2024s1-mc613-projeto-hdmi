module spriteObjeto1 (
	input clk,
	input reset,
	input [9:0] x, y, sprite_x, sprite_y,
	input vsync,
	output reg color,
	output reg drawing
);

parameter [6:0] sprite_width = (16*9) + (4*8);  //172
parameter  sprite_height = 16;
reg [0:sprite_width-1] bmap [sprite_height];
initial begin
	bmap[0]  = 172'b1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_0_0_0_0_0_0_0_0_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_0_0_0_0;
	bmap[1]  = 172'b1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_0_0_0_0_0_0_0_0_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_0_0_0_0;
	bmap[2]  = 172'b1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_0_0_0_0_0_0_0_0_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1;
	bmap[3]  = 172'b1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_0_0_0_0_0_0_0_0_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1;
	bmap[4]  = 172'b1_1_1_1_0_0_0_0_0_0_0_0_0_0_0_0__0000__1_1_1_1_0_0_0_0_0_0_0_0_1_1_1_1__0000__1_1_1_1_0_0_1_1_1_1_0_0_1_1_1_1__0000__1_1_1_1_0_0_0_0_0_0_0_0_0_0_0_0__0000__1_1_1_1_0_0_0_0_0_0_0_0_1_1_1_1__0000__0_1_1_1_1_0_0_0_0_0_0_0_1_1_1_0__0000__1_1_1_1_0_0_0_0_0_0_0_0_0_0_0_0__0000__1_1_1_1_0_0_0_0_0_0_0_0_1_1_1_1;
	bmap[5]  = 172'b1_1_1_1_0_0_0_0_0_0_0_0_0_0_0_0__0000__1_1_1_1_0_0_0_0_0_0_0_0_1_1_1_1__0000__1_1_1_1_0_0_1_1_1_1_0_0_1_1_1_1__0000__1_1_1_1_0_0_0_0_0_0_0_0_0_0_0_0__0000__1_1_1_1_0_0_0_0_0_0_0_0_1_1_1_1__0000__0_1_1_1_1_0_0_0_0_0_0_1_1_1_1_0__0000__1_1_1_1_0_0_0_0_0_0_0_0_0_0_0_0__0000__1_1_1_1_0_0_0_0_0_0_0_0_1_1_1_1;
	bmap[6]  = 172'b1_1_1_1_0_0_0_0_0_0_0_0_0_0_0_0__0000__1_1_1_1_0_0_0_0_0_0_0_0_1_1_1_1__0000__1_1_1_1_0_0_1_1_1_1_0_0_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_0_0_0_0_0_0_0_0_1_1_1_1__0000__0_0_1_1_1_1_0_0_0_0_1_1_1_1_0_0__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_0_0_0_0_0_0_0_0_1_1_1_1;
	bmap[7]  = 172'b1_1_1_1_0_0_0_0_0_0_0_0_0_0_0_0__0000__1_1_1_1_0_0_0_0_0_0_0_0_1_1_1_1__0000__1_1_1_1_0_0_1_1_1_1_0_0_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_0_0_0_0_0_0_0_0_1_1_1_1__0000__0_0_1_1_1_1_0_0_0_0_1_1_1_1_0_0__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_0_0_0_0_0_0_0_0_1_1_1_1;
	bmap[8]  = 172'b1_1_1_1_0_0_0_0_0_0_1_1_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_0_0_1_1_1_1_0_0_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_0_0_0_0_0_0_0_0_1_1_1_1__0000__0_0_0_1_1_1_1_0_0_1_1_1_1_0_0_0__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1;
	bmap[9]  = 172'b1_1_1_1_0_0_0_0_0_0_1_1_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_0_0_1_1_1_1_0_0_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_0_0_0_0_0_0_0_0_1_1_1_1__0000__0_0_0_1_1_1_1_0_0_1_1_1_1_0_0_0__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1;
	bmap[10] = 172'b1_1_1_1_0_0_0_0_0_0_0_0_1_1_1_1__0000__1_1_1_1_0_0_0_0_0_0_0_0_1_1_1_1__0000__1_1_1_1_0_0_1_1_1_1_0_0_1_1_1_1__0000__1_1_1_1_0_0_0_0_0_0_0_0_0_0_0_0__0000__1_1_1_1_0_0_0_0_0_0_0_0_1_1_1_1__0000__0_0_0_0_1_1_1_1_1_1_1_1_0_0_0_0__0000__1_1_1_1_0_0_0_0_0_0_0_0_0_0_0_0__0000__1_1_1_1_1_1_1_1_1_1_1_1_0_0_0_0;
	bmap[11] = 172'b1_1_1_1_0_0_0_0_0_0_0_0_1_1_1_1__0000__1_1_1_1_0_0_0_0_0_0_0_0_1_1_1_1__0000__1_1_1_1_0_0_1_1_1_1_0_0_1_1_1_1__0000__1_1_1_1_0_0_0_0_0_0_0_0_0_0_0_0__0000__1_1_1_1_0_0_0_0_0_0_0_0_1_1_1_1__0000__0_0_0_0_1_1_1_1_1_1_1_1_0_0_0_0__0000__1_1_1_1_0_0_0_0_0_0_0_0_0_0_0_0__0000__1_1_1_1_1_1_1_1_1_1_1_1_0_0_0_0;
	bmap[12] = 172'b1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_0_0_0_0_0_0_0_0_1_1_1_1__0000__1_1_1_1_0_0_1_1_1_1_0_0_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__0_0_0_0_0_1_1_1_1_1_1_0_0_0_0_0__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_0_0_0_0_1_1_1_1_0_0_0_0;
	bmap[13] = 172'b1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_0_0_0_0_0_0_0_0_1_1_1_1__0000__1_1_1_1_0_0_1_1_1_1_0_0_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__0_0_0_0_0_1_1_1_1_1_1_0_0_0_0_0__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_0_0_0_0_0_1_1_1_1_1_0_0;
	bmap[14] = 172'b1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_0_0_0_0_0_0_0_0_1_1_1_1__0000__1_1_1_1_0_0_1_1_1_1_0_0_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__0_0_0_0_0_0_1_1_1_1_0_0_0_0_0_0__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_0_0_0_0_0_0_1_1_1_1_1_0;
	bmap[15] = 172'b1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_0_0_0_0_0_0_0_0_1_1_1_1__0000__1_1_1_1_0_0_1_1_1_1_0_0_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__0_0_0_0_0_0_1_1_1_1_0_0_0_0_0_0__0000__1_1_1_1_1_1_1_1_1_1_1_1_1_1_1_1__0000__1_1_1_1_0_0_0_0_0_0_0_0_1_1_1_1;
end

reg [$clog2(sprite_width)-1:0] bmap_x;
reg [$clog2(sprite_height)-1:0] bmap_y;

reg [9:0] sprite_x_reg, sprite_y_reg;
always @ (negedge vsync) begin
	sprite_x_reg = sprite_x;
	sprite_y_reg = sprite_y;
end 

reg sprite_active_y, sprite_active_x, sprite_end, line_end;

always @ (x, y) begin
	sprite_active_y = (y >= sprite_y_reg) && (y < sprite_y_reg + sprite_height);
	sprite_active_x = (x >= sprite_x_reg) && (x < sprite_x_reg + sprite_width);
	bmap_x = x - sprite_x_reg;
	bmap_y = y - sprite_y_reg;
	drawing = (sprite_active_y && sprite_active_x) ? 1 : 0;
	color = (sprite_active_y && sprite_active_x) ? bmap[bmap_y][bmap_x] : 0;
end

endmodule